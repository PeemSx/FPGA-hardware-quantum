module hadamard(
    input clk,
    input reset,
    
);


endmodule